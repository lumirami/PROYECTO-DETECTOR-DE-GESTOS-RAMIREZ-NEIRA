doscientos_inst : doscientos PORT MAP (
		result	 => result_sig
	);
